io_in_inst : io_in PORT MAP (
		datain	 => datain_sig,
		inclock	 => inclock_sig,
		inclocken	 => inclocken_sig,
		dataout_h	 => dataout_h_sig,
		dataout_l	 => dataout_l_sig
	);
